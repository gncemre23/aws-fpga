
//TODO draw new diagram regarding the new code
/* ================== Heavy hash block ================================= */
/*           Block_header            Matrix               Target         */
/*                |                     |                    |           */
/*                |                     |                    |           */
/*                |                     |                    |           */
/*       +--------+---------------------+--------------------+---------+ */
/*       |        |                     v                    |         | */
/*       |        v                +----------+              v         | */
/* start |   +----------+          |          |        +-----------+   | */
/* ------+-->| nonce_gen+--------->|heavy_hash+------->|comparator |   | */
/*       |   +----+-----+          |          |        +-----+-----+   | */
/*       |                         +----------+              |         | */
/*       |                               |                   |         | */
/*       +--------+----------------------|-------------------+---------+ */
/*                                       |                   |           */
/*                                       |                   |           */
/*                                       v                   v           */
/*                                     nonce               result        */
/* ================== Heavy hash block ================================= */
`timescale  1ns / 1ps
module heavy_hash_blk
  #(
     parameter NONCE_COEF = 1,
     parameter WCOUNT = 4
   )
   (
     //!global clk
     input logic clk,
     //!global reset
     input logic rst,

     //! start signal for new block operations
     input logic start,

     //! stop signal
     input logic stop,

     //! 32-bit block header input (dout data from block_header fifo)
     input logic [31:0] block_header,

     //! 32-bit matrix_in input from matrix_fifo
     input logic [31:0] matrix_in,

     //! 32-bit target input
     input logic [31:0] target,

     //! 32-bit size calculated by software
     input logic [31:0] nonce_size,

     //! matrix fifo write enable
     input logic matrix_we,

     //! nonce output generated by nonce_gen
     output logic [31:0] nonce,

     //! result stating if the output of heavy hash is less than the target
     //! 1 : less than target (objective)
     //! 0 : greater than target
     output logic result,

     //! acknowledge signal stating ready to recieve start signal
     output logic stop_ack,

     //! status
     output logic [1:0] status,

     output logic [255:0] hash_out,
     output logic hash_out_we

   );


  //internal signals
  logic hashin_fifo_in_we;
  logic [63:0] hashin_fifo_in_din;
  logic hashin_fifo_in_full;
  logic matrix_fifo_in_full;
  logic hashout_fifo_re;
  logic [255:0] hashout_fifo_out_dout;
  logic hash_out_empty;
  logic nonce_fifo_we;
  logic nonce_fifo_full;
  logic stop_ack_comp;
  logic stop_ack_nonce;
  logic [31:0] nonce_fifo_din;
  logic [255:0] zero_reg  = 256'd0;
  logic heavy_hash_all_empty;
  logic [31:0] nonce_end;


  assign stop_ack = stop_ack_comp & stop_ack_nonce;

  assign hash_out_we = hashout_fifo_re;

  always_comb begin : blockName
    if(result)
      status = 1;
    else if(nonce < nonce_end)
      status = 0;
    else
      status = 2;
  end

  nonce_gen
    #(
      .NONCE_COEF ( NONCE_COEF )
    )
    nonce_gen_dut (
      .clk (clk ),
      .rst (rst ),
      .start (start ),
      .stop (stop ),
      .block_header (block_header ),
      .nonce_size (nonce_size ),
      .hashin_fifo_in_we (hashin_fifo_in_we ),
      .hashin_fifo_in_din (hashin_fifo_in_din ),
      .hashin_fifo_in_full (hashin_fifo_in_full ),
      .nonce_fifo_full (nonce_fifo_full ),
      .nonce_fifo_din (nonce_fifo_din ),
      .nonce_fifo_we (nonce_fifo_we ),
      .stop_ack_nonce  ( stop_ack_nonce),
      .nonce_end(nonce_end)
    );


  heavy_hash
    #(
      .WCOUNT ( WCOUNT )
    )
    heavy_hash_dut (
      .clk (clk ),
      .rst (rst ),
      .hashin_fifo_in_we (hashin_fifo_in_we ),
      .hashin_fifo_in_din (hashin_fifo_in_din ),
      .hashin_fifo_in_full (hashin_fifo_in_full ),
      .matrix_fifo_in_we (matrix_we ),
      .matrix_fifo_in_din (matrix_in ),
      // not expecting to be full. TODO: matrix fifo will be taken out from heavy hash
      // only one fifo is enough
      .matrix_fifo_in_full (matrix_fifo_in_full ),
      .hashout_fifo_out_re (hashout_fifo_re ),
      .hashout_fifo_out_dout (hash_out ),
      .hashout_fifo_out_empty  ( hash_out_empty),
      .nonce_fifo_din(nonce_fifo_din),
      .nonce_fifo_we(nonce_fifo_we),
      .nonce_fifo_full(nonce_fifo_full),
      .nonce(nonce),
      .heavy_hash_all_empty(heavy_hash_all_empty)
    );

  comparator
    comparator_inst(
      .clk (clk ),
      .rst (rst ),
      .target (target ),
      .start (start ),
      .stop(stop ),
      .stop_ack_comp (stop_ack_comp ),
      .heavy_hash_all_empty (heavy_hash_all_empty ),
      .hashout_fifo_re (hashout_fifo_re ),
      .hash_out (hash_out ),
      .hash_out_empty (hash_out_empty ),
      .result  ( result)
    );





endmodule
